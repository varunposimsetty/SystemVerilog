module traffic (
    
);
    
endmodule